LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fastSram is 
	port(
		
	)
	
	
	
architecture bhv of fastSram is
begin

end bhv;