LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fileSystem is
	port(
		
	);
end fileSystem;

architecture bhv of fileSystem is
begin
	
end bhv;